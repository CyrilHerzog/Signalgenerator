
/*
    Module  : BARREL_SHIFTER_DEFINES
    Version : 1.1
    Author  : Herzog Cyril
    Date    : 09.11.2024

*/


`ifndef BARREL_SHIFTER_DEFINES_VH
`define BARREL_SHIFTER_DEFINES_VH


`define SHIFT_MODE_BIDIRECTIONAL 0
`define SHIFT_MODE_RIGHT         1
`define SHIFT_MODE_LEFT          2


`endif /* BARREL_SHIFTER_DEFINES */
